module regn ( 
	d,
	clk,
	rin,
	q
	) ;

input [1:0] d;
input  clk;
input  rin;
inout [1:0] q;
