module control_registers ( 
	t,
	i,
	x,
	y,
	rin,
	rout
	) ;

input [3:0] t;
input [3:0] i;
input [2:0] x;
input [2:0] y;
inout [2:0] rin;
inout [2:0] rout;
