module control_alu ( 
	t,
	i,
	ain,
	gin,
	gout,
	addsub
	) ;

input [3:0] t;
input [3:0] i;
inout  ain;
inout  gin;
inout  gout;
inout  addsub;
