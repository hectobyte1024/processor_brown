module gal2_register_decoder ( 
	rx_in,
	ry_in,
	x,
	y
	) ;

input [1:0] rx_in;
input [1:0] ry_in;
inout [2:0] x;
inout [2:0] y;
